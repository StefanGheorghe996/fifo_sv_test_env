library verilog;
use verilog.vl_types.all;
entity fifo_generator is
end fifo_generator;
