library verilog;
use verilog.vl_types.all;
entity fifo_packet_sv_unit is
end fifo_packet_sv_unit;
