library verilog;
use verilog.vl_types.all;
entity fifo_include_sv_unit is
end fifo_include_sv_unit;
