library verilog;
use verilog.vl_types.all;
entity fifo_generator_sv_unit is
end fifo_generator_sv_unit;
