package fifo_include;
`include "env/fifo_if.sv"
`include "env/fifo_base_unit.sv"
`include "env/fifo_packet.sv"
`include "env/fifo_driver.sv"
`include "env/fifo_generator.sv"
`include "env/fifo_tb.sv"
`include "env/fifo_environment.sv"
endpackage