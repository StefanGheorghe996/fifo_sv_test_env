library verilog;
use verilog.vl_types.all;
entity fifo_test_basic_sv_unit is
end fifo_test_basic_sv_unit;
