library verilog;
use verilog.vl_types.all;
entity fifo_driver is
end fifo_driver;
