library verilog;
use verilog.vl_types.all;
entity fifo_base_unit_sv_unit is
end fifo_base_unit_sv_unit;
