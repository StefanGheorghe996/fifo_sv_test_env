library verilog;
use verilog.vl_types.all;
entity fifo_tb_sv_unit is
end fifo_tb_sv_unit;
