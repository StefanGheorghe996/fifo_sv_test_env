library verilog;
use verilog.vl_types.all;
entity fifo_driver_sv_unit is
end fifo_driver_sv_unit;
